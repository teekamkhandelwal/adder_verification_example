//transection
class transaction;
  rand bit [3:0]a,b;
  bit [4:0] sum;
endclass
